`timescale 1ns / 1ps

module top(
    //input
	kasia
    //output
	
    );
    
    
endmodule
